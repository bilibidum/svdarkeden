/home/darkeden/vs/bin
