/home/rafael/darkeden/vs/bin
